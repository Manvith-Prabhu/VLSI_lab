* NMOS Resistive Load Inverter

.include ./t14y_tsmc_025_level3.txt

m1 vout vin 0 0 cmosn l=0.5u w=10u
r1 vdd vout 10000

v_dd vdd 0 5
v_in vin 0 PULSE(0 5 0 0.0001n 0.0001n 10m 20m)


.control
    dc v_in 0 5 0.01
    
    **** FOR WIDTH MANIPULATION
    *foreach wid 1e-7 1e-5 1e-4
    *alter m1 w = $wen
    *run
    *end
    ***********************
    
    foreach len 1e-7 1e-5 1e-4
    alter m1 l = $len
    run
    end
    
    foreach iter 1 2 3 
    setplot dc$iter
    plot vout
    plot -v_dd#branch
    plot deriv(vout)
    end
.endc

.end





