magic
tech scmos
timestamp 1699718400
<< polysilicon >>
rect 7 19 9 21
rect 7 3 9 13
rect 7 -2 9 0
<< ndiffusion >>
rect 4 0 7 3
rect 9 0 11 3
rect 15 0 16 3
<< pdiffusion >>
rect 4 16 7 19
rect 0 13 7 16
rect 9 17 16 19
rect 9 13 11 17
rect 15 13 16 17
<< metal1 >>
rect 0 24 7 27
rect 11 24 17 27
rect 0 20 4 24
rect 11 3 15 13
rect 0 -4 4 -1
rect 0 -5 16 -4
rect 0 -7 6 -5
rect 10 -7 16 -5
<< ntransistor >>
rect 7 0 9 3
<< ptransistor >>
rect 7 13 9 19
<< polycontact >>
rect 3 7 7 11
<< ndcontact >>
rect 0 -1 4 3
rect 11 -1 15 3
<< pdcontact >>
rect 0 16 4 20
rect 11 13 15 17
<< psubstratepcontact >>
rect 6 -9 10 -5
<< nsubstratencontact >>
rect 7 24 11 28
<< labels >>
rlabel metal1 11 7 15 11 7 out
rlabel polycontact 3 7 7 11 3 in
rlabel nsubstratencontact 7 24 11 28 5 vdd
rlabel psubstratepcontact 6 -9 10 -5 1 vss
<< end >>
