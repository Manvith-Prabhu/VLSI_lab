* SPICE3 file created from nor2.ext - technology: scmos
.include ./t14y_tsmc_025_level3.txt
.option scale=1u

M1000 a_7_18# A Vdd Vdd cmosp w=6 l=2
+  ad=54 pd=30 as=32 ps=24
M1001 Vout B a_7_18# Vdd cmosp w=6 l=2
+  ad=36 pd=26 as=0 ps=0
M1002 Vout A Gnd Gnd cmosn w=3 l=2
+  ad=31 pd=26 as=44 ps=40
M1003 Gnd B Vout Gnd cmosn w=3 l=2
+  ad=0 pd=0 as=0 ps=0
C0 Gnd Gnd 4.32fF
C1 Vout Gnd 4.65fF
C2 B Gnd 7.07fF
C3 A Gnd 7.07fF
C4 Vdd Gnd 3.43fF


vdd Vdd 0 5
gnd Gnd 0 0
va A 0 PULSE(0 5 0 0 0 4n 8n)
vb B 0 PULSE(0 5 0 0 0 2n 4n)

.control
tran 0.01p 10n
setplot tran
plot A B Vout

.endc

.end
 
