* SPICE3 file created from nor3.ext - technology: scmos

.option scale=1u

M1000 a_7_18# A Vdd Vdd pfet w=6 l=2
+  ad=54 pd=30 as=32 ps=24
M1001 a_18_18# B a_7_18# Vdd pfet w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1002 Vout C a_18_18# Vdd pfet w=6 l=2
+  ad=36 pd=26 as=0 ps=0
M1003 Vout A gnd Gnd nfet w=3 l=2
+  ad=59 pd=50 as=44 ps=40
M1004 gnd B Vout Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 Vout C gnd Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
C0 gnd Gnd 4.18fF
C1 Vout Gnd 6.44fF
C2 C Gnd 7.07fF
C3 B Gnd 7.07fF
C4 A Gnd 7.07fF
C5 Vdd Gnd 3.43fF
